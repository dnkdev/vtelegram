module media
